//////////////////////////////////////////////////////////////////////////
//                                                                      //
//   Modulename :  ex_stage.v                                           //
//                                                                      //
//  Description :  instruction execute (EX) stage of the pipeline;      //
//                 given the instruction command code CMD, select the   //
//                 proper input A and B for the ALU, compute the result,// 
//                 and compute the condition for branches, and pass all //
//                 the results down the pipeline. MWB                   // 
//                                                                      //
//                                                                      //
//////////////////////////////////////////////////////////////////////////
`ifndef __ALU_FU_V__
`define __ALU_FU_V__

//`timescale 1ns/100ps

//
// The ALU
//
// given the command code CMD and proper operands A and B, compute the
// result of the instruction
//
// This module is purely combinational
//
module alu(
	input [`XLEN-1:0] opa,
	input [`XLEN-1:0] opb,
	ALU_FUNC     func,

	output logic [`XLEN-1:0] result
);
	wire signed [`XLEN-1:0] signed_opa, signed_opb;
	// wire signed [2*`XLEN-1:0] signed_mul, mixed_mul;
	// wire        [2*`XLEN-1:0] unsigned_mul;
	assign signed_opa = opa;
	assign signed_opb = opb;
	// assign signed_mul = signed_opa * signed_opb;
	// assign unsigned_mul = opa * opb;
	// assign mixed_mul = signed_opa * opb;

	always_comb begin
		case (func)
			ALU_ADD:      result = opa + opb;
			ALU_SUB:      result = opa - opb;
			ALU_AND:      result = opa & opb;
			ALU_SLT:      result = signed_opa < signed_opb;
			ALU_SLTU:     result = opa < opb;
			ALU_OR:       result = opa | opb;
			ALU_XOR:      result = opa ^ opb;
			ALU_SRL:      result = opa >> opb[4:0];
			ALU_SLL:      result = opa << opb[4:0];
			ALU_SRA:      result = signed_opa >>> opb[4:0]; // arithmetic from logical shift
			// ALU_MUL:      result = signed_mul[`XLEN-1:0];
			// ALU_MULH:     result = signed_mul[2*`XLEN-1:`XLEN];
			// ALU_MULHSU:   result = mixed_mul[2*`XLEN-1:`XLEN];
			// ALU_MULHU:    result = unsigned_mul[2*`XLEN-1:`XLEN];

			default:      result = `XLEN'hfacebeec;  // here to prevent latches
		endcase
	end
endmodule // alu

//
// BrCond module
//
// Given the instruction code, compute the proper condition for the
// instruction; for branches this condition will indicate whether the
// target is taken.
//
// This module is purely combinational
//
module brcond(// Inputs
	input [`XLEN-1:0] rs1,    // Value to check against condition
	input [`XLEN-1:0] rs2,
	input  [2:0] func,  // Specifies which condition to check

	output logic cond    // 0/1 condition result (False/True)
);

	logic signed [`XLEN-1:0] signed_rs1, signed_rs2;
	assign signed_rs1 = rs1;
	assign signed_rs2 = rs2;
	always_comb begin
		cond = 0;
		case (func)
			3'b000: cond = signed_rs1 == signed_rs2;  // BEQ
			3'b001: cond = signed_rs1 != signed_rs2;  // BNE
			3'b100: cond = signed_rs1 < signed_rs2;   // BLT
			3'b101: cond = signed_rs1 >= signed_rs2;  // BGE
			3'b110: cond = rs1 < rs2;                 // BLTU
			3'b111: cond = rs1 >= rs2;                // BGEU
		endcase
	end
	
endmodule // brcond


module alu_fu(
	input clock,               // system clock
	input reset,               // system reset
	input enable,
	input squash_in,
	input IS_EX_PACKET   is_ex_packet_in,
	output EX_BP_PACKET  ex_bp_packet_out,
	output EX_CP_PACKET  ex_cp_packet
);
	EX_CP_PACKET  ex_packet_out;
	EX_BP_PACKET  ex_bp_packet;
	logic [`XLEN-1:0] alu_result;
	// Pass-throughs
    assign ex_packet_out.inst = is_ex_packet_in.inst;
	assign ex_packet_out.dest_reg_idx = is_ex_packet_in.dest_reg_idx;
	assign ex_packet_out.halt = is_ex_packet_in.halt;
	assign ex_packet_out.illegal = is_ex_packet_in.illegal;
	assign ex_packet_out.valid = is_ex_packet_in.valid;
	assign ex_packet_out.done = is_ex_packet_in.valid;
    assign ex_packet_out.Tag = is_ex_packet_in.Tag;

	

	// assign ex_packet_out.mem_size = is_ex_packet_in.inst.r.funct3;

	logic [`XLEN-1:0] opa_mux_out, opb_mux_out;
	logic brcond_result;
	//
	// ALU opA mux
	//
	always_comb begin
		opa_mux_out = `XLEN'hdeadfbac;
		case (is_ex_packet_in.opa_select)
			OPA_IS_RS1:  opa_mux_out = is_ex_packet_in.rs1_value;
			OPA_IS_NPC:  opa_mux_out = is_ex_packet_in.NPC;
			OPA_IS_PC:   opa_mux_out = is_ex_packet_in.PC;
			OPA_IS_ZERO: opa_mux_out = 0;
		endcase
	end

	 //
	 // ALU opB mux
	 //
	always_comb begin
		// Default value, Set only because the case isnt full.  If you see this
		// value on the output of the mux you have an invalid opb_select
		opb_mux_out = `XLEN'hfacefeed;
		case (is_ex_packet_in.opb_select)
			OPB_IS_RS2:   opb_mux_out = is_ex_packet_in.rs2_value;
			OPB_IS_I_IMM: opb_mux_out = `RV32_signext_Iimm(is_ex_packet_in.inst);
			OPB_IS_S_IMM: opb_mux_out = `RV32_signext_Simm(is_ex_packet_in.inst);
			OPB_IS_B_IMM: opb_mux_out = `RV32_signext_Bimm(is_ex_packet_in.inst);
			OPB_IS_U_IMM: opb_mux_out = `RV32_signext_Uimm(is_ex_packet_in.inst);
			OPB_IS_J_IMM: opb_mux_out = `RV32_signext_Jimm(is_ex_packet_in.inst);
		endcase 
	end

	//
	// instantiate the ALU
	//
	alu alu_0 (// Inputs
		.opa(opa_mux_out),
		.opb(opb_mux_out),
		.func(is_ex_packet_in.alu_func),

		// Output
		.result(alu_result)
	);

	 //
	 // instantiate the branch condition tester
	 //
	brcond brcond (// Inputs
		.rs1(is_ex_packet_in.rs1_value), 
		.rs2(is_ex_packet_in.rs2_value),
		.func(is_ex_packet_in.inst.b.funct3), // inst bits to determine check

		// Output
		.cond(brcond_result)
	);

	// mux to select writeback data
	assign ex_packet_out.Value = is_ex_packet_in.uncond_branch
		                          | (is_ex_packet_in.cond_branch & brcond_result) ? is_ex_packet_in.PC + 4 : alu_result;

	//mux to select next PC
	assign ex_packet_out.NPC = is_ex_packet_in.uncond_branch
		                          | (is_ex_packet_in.cond_branch & brcond_result) ? alu_result : is_ex_packet_in.PC + 4;

	 // ultimate "take branch" signal:
	 //	unconditional, or conditional and the condition is true
	assign ex_packet_out.take_branch = (ex_packet_out.NPC != is_ex_packet_in.NPC) & ex_bp_packet.br_en;

	// go to BP
	assign ex_bp_packet.PC = is_ex_packet_in.PC;
	assign ex_bp_packet.br_en = is_ex_packet_in.uncond_branch
	               				| is_ex_packet_in.cond_branch;
	assign ex_bp_packet.con_br_en = is_ex_packet_in.cond_branch;
	assign ex_bp_packet.con_br_taken = is_ex_packet_in.cond_branch & brcond_result;
    assign ex_bp_packet.tg_pc = alu_result;

	// synopsys sync_set_reset "reset"
	always_ff @(posedge clock) begin
		if (reset)begin
			ex_cp_packet.Value <= `SD 0;
			ex_cp_packet.NPC <= `SD 0;
			ex_cp_packet.take_branch <= `SD 0;
			ex_cp_packet.inst <= `SD `NOP;
			ex_cp_packet.dest_reg_idx <= `SD `ZERO_REG;
			ex_cp_packet.halt <= `SD `FALSE;
			ex_cp_packet.illegal <= `SD `FALSE;
			ex_cp_packet.valid <= `SD 0;
			ex_cp_packet.done <= `SD 0;
			ex_cp_packet.Tag <= `SD 0;
		end
		else if (squash_in) begin
			ex_cp_packet.Value <= `SD 0;
			ex_cp_packet.NPC <= `SD 0;
			ex_cp_packet.take_branch <= `SD 0;
			ex_cp_packet.inst <= `SD `NOP;
			ex_cp_packet.dest_reg_idx <= `SD `ZERO_REG;
			ex_cp_packet.halt <= `SD `FALSE;
			ex_cp_packet.illegal <= `SD `FALSE;
			ex_cp_packet.valid <= `SD 0;
			ex_cp_packet.done <= `SD 0;
			ex_cp_packet.Tag <= `SD 0;
		end
		else if (enable) begin
			ex_cp_packet <= `SD ex_packet_out;
		end
	end

	// synopsys sync_set_reset "reset"
	always_ff @(posedge clock) begin
		if (reset) begin
			ex_bp_packet_out <= `SD 0;
		end
		else if (squash_in) begin
			ex_bp_packet_out <= `SD 0;
		end
		else if (enable) begin
			ex_bp_packet_out <= `SD ex_bp_packet;
		end
		else begin
			ex_bp_packet_out <= `SD 0;
		end
	end

endmodule // module ex_stage
`endif // __ALU_FU_V__
